module MatissaAdder48(input wire[55:8]  A,B,
                      input wire        ct,
                      output wire[55:8] out);

    wire[28:0] h0a,h0b,h1a,h1b;
    wire[31:0] thout;
    

endmodule