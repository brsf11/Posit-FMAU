module MatissaWallaceTree28x28();

endmodule