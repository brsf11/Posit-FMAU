module Compressor73(input wire  x1,x2,x3,x4,x5,x6,x7,
                    output reg s,c1,c2);

endmodule