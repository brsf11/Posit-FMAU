module UnsignedMultiplier7x7(input wire[6:0]   A,B,
                             output wire[13:0] out);

endmodule