module MatissaWallaceTree28x28(input wire[13:0]  PP11,
                               input wire[20:7]  PP12,PP21,
                               input wire[27:14] PP13,PP22,PP31,
                               input wire[34:21] PP14,PP23,PP32,PP41,
                               input wire[41:28] PP24,PP33,PP42,
                               input wire[48:35] PP34,PP43,
                               input wire[55:42] PP44,
                               input wire[1:0]   op,
                               output wire[55:0] out);

    

endmodule