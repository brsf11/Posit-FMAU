module Compressor73(input wire  x1,x2,x3,x4,x5,x6,x7,
                    output reg  s,c1,c2);

    always @(*) begin
        case({x1,x2,x3,x4,x5,x6,x7})
            7'b0000000: {c1,c2,s} = 3'b000;
            7'b0000001: {c1,c2,s} = 3'b001;
            7'b0000010: {c1,c2,s} = 3'b001;
            7'b0000011: {c1,c2,s} = 3'b010;
            7'b0000100: {c1,c2,s} = 3'b001;
            7'b0000101: {c1,c2,s} = 3'b010;
            7'b0000110: {c1,c2,s} = 3'b010;
            7'b0000111: {c1,c2,s} = 3'b011;
            7'b0001000: {c1,c2,s} = 3'b001;
            7'b0001001: {c1,c2,s} = 3'b010;
            7'b0001010: {c1,c2,s} = 3'b010;
            7'b0001011: {c1,c2,s} = 3'b011;
            7'b0001100: {c1,c2,s} = 3'b010;
            7'b0001101: {c1,c2,s} = 3'b011;
            7'b0001110: {c1,c2,s} = 3'b011;
            7'b0001111: {c1,c2,s} = 3'b100;
            7'b0010000: {c1,c2,s} = 3'b001;
            7'b0010001: {c1,c2,s} = 3'b010;
            7'b0010010: {c1,c2,s} = 3'b010;
            7'b0010011: {c1,c2,s} = 3'b011;
            7'b0010100: {c1,c2,s} = 3'b010;
            7'b0010101: {c1,c2,s} = 3'b011;
            7'b0010110: {c1,c2,s} = 3'b011;
            7'b0010111: {c1,c2,s} = 3'b100;
            7'b0011000: {c1,c2,s} = 3'b010;
            7'b0011001: {c1,c2,s} = 3'b011;
            7'b0011010: {c1,c2,s} = 3'b011;
            7'b0011011: {c1,c2,s} = 3'b100;
            7'b0011100: {c1,c2,s} = 3'b011;
            7'b0011101: {c1,c2,s} = 3'b100;
            7'b0011110: {c1,c2,s} = 3'b100;
            7'b0011111: {c1,c2,s} = 3'b101;

            7'b0100000: {c1,c2,s} = 3'b001;
            7'b0100001: {c1,c2,s} = 3'b010;
            7'b0100010: {c1,c2,s} = 3'b010;
            7'b0100011: {c1,c2,s} = 3'b011;
            7'b0100100: {c1,c2,s} = 3'b010;
            7'b0100101: {c1,c2,s} = 3'b011;
            7'b0100110: {c1,c2,s} = 3'b011;
            7'b0100111: {c1,c2,s} = 3'b100;
            7'b0101000: {c1,c2,s} = 3'b010;
            7'b0101001: {c1,c2,s} = 3'b011;
            7'b0101010: {c1,c2,s} = 3'b011;
            7'b0101011: {c1,c2,s} = 3'b100;
            7'b0101100: {c1,c2,s} = 3'b011;
            7'b0101101: {c1,c2,s} = 3'b100;
            7'b0101110: {c1,c2,s} = 3'b100;
            7'b0101111: {c1,c2,s} = 3'b101;
            7'b0110000: {c1,c2,s} = 3'b010;
            7'b0110001: {c1,c2,s} = 3'b011;
            7'b0110010: {c1,c2,s} = 3'b011;
            7'b0110011: {c1,c2,s} = 3'b100;
            7'b0110100: {c1,c2,s} = 3'b011;
            7'b0110101: {c1,c2,s} = 3'b100;
            7'b0110110: {c1,c2,s} = 3'b100;
            7'b0110111: {c1,c2,s} = 3'b101;
            7'b0111000: {c1,c2,s} = 3'b011;
            7'b0111001: {c1,c2,s} = 3'b100;
            7'b0111010: {c1,c2,s} = 3'b100;
            7'b0111011: {c1,c2,s} = 3'b101;
            7'b0111100: {c1,c2,s} = 3'b100;
            7'b0111101: {c1,c2,s} = 3'b101;
            7'b0111110: {c1,c2,s} = 3'b101;
            7'b0111111: {c1,c2,s} = 3'b110;

            7'b1000000: {c1,c2,s} = 3'b001;
            7'b1000001: {c1,c2,s} = 3'b010;
            7'b1000010: {c1,c2,s} = 3'b010;
            7'b1000011: {c1,c2,s} = 3'b011;
            7'b1000100: {c1,c2,s} = 3'b010;
            7'b1000101: {c1,c2,s} = 3'b011;
            7'b1000110: {c1,c2,s} = 3'b011;
            7'b1000111: {c1,c2,s} = 3'b100;
            7'b1001000: {c1,c2,s} = 3'b010;
            7'b1001001: {c1,c2,s} = 3'b011;
            7'b1001010: {c1,c2,s} = 3'b011;
            7'b1001011: {c1,c2,s} = 3'b100;
            7'b1001100: {c1,c2,s} = 3'b011;
            7'b1001101: {c1,c2,s} = 3'b100;
            7'b1001110: {c1,c2,s} = 3'b100;
            7'b1001111: {c1,c2,s} = 3'b101;
            7'b1010000: {c1,c2,s} = 3'b010;
            7'b1010001: {c1,c2,s} = 3'b011;
            7'b1010010: {c1,c2,s} = 3'b011;
            7'b1010011: {c1,c2,s} = 3'b100;
            7'b1010100: {c1,c2,s} = 3'b011;
            7'b1010101: {c1,c2,s} = 3'b100;
            7'b1010110: {c1,c2,s} = 3'b100;
            7'b1010111: {c1,c2,s} = 3'b101;
            7'b1011000: {c1,c2,s} = 3'b011;
            7'b1011001: {c1,c2,s} = 3'b100;
            7'b1011010: {c1,c2,s} = 3'b100;
            7'b1011011: {c1,c2,s} = 3'b101;
            7'b1011100: {c1,c2,s} = 3'b100;
            7'b1011101: {c1,c2,s} = 3'b101;
            7'b1011110: {c1,c2,s} = 3'b101;
            7'b1011111: {c1,c2,s} = 3'b110;

            7'b1100000: {c1,c2,s} = 3'b010;
            7'b1100001: {c1,c2,s} = 3'b011;
            7'b1100010: {c1,c2,s} = 3'b011;
            7'b1100011: {c1,c2,s} = 3'b100;
            7'b1100100: {c1,c2,s} = 3'b011;
            7'b1100101: {c1,c2,s} = 3'b100;
            7'b1100110: {c1,c2,s} = 3'b100;
            7'b1100111: {c1,c2,s} = 3'b101;
            7'b1101000: {c1,c2,s} = 3'b011;
            7'b1101001: {c1,c2,s} = 3'b100;
            7'b1101010: {c1,c2,s} = 3'b100;
            7'b1101011: {c1,c2,s} = 3'b101;
            7'b1101100: {c1,c2,s} = 3'b100;
            7'b1101101: {c1,c2,s} = 3'b101;
            7'b1101110: {c1,c2,s} = 3'b101;
            7'b1101111: {c1,c2,s} = 3'b110;
            7'b1110000: {c1,c2,s} = 3'b011;
            7'b1110001: {c1,c2,s} = 3'b100;
            7'b1110010: {c1,c2,s} = 3'b100;
            7'b1110011: {c1,c2,s} = 3'b101;
            7'b1110100: {c1,c2,s} = 3'b100;
            7'b1110101: {c1,c2,s} = 3'b101;
            7'b1110110: {c1,c2,s} = 3'b101;
            7'b1110111: {c1,c2,s} = 3'b110;
            7'b1111000: {c1,c2,s} = 3'b100;
            7'b1111001: {c1,c2,s} = 3'b101;
            7'b1111010: {c1,c2,s} = 3'b101;
            7'b1111011: {c1,c2,s} = 3'b110;
            7'b1111100: {c1,c2,s} = 3'b101;
            7'b1111101: {c1,c2,s} = 3'b110;
            7'b1111110: {c1,c2,s} = 3'b110;
            7'b1111111: {c1,c2,s} = 3'b111;
            default:    {c1,c2,s} = 3'b000;
        endcase
    end

endmodule