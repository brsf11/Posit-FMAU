module UnsignedMultiplier7x7();

endmodule