module WallaceTreeSigned8x8(input wire[11:0] pp00,pp03,
                            input wire[12:0] pp01,pp02);

    wire
    
endmodule